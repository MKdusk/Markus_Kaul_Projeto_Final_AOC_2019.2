LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SomadorPC IS
PORT(
	   AddIn : in STD_LOGIC_VECTOR(7 DOWNTO 0);
		AddInTwo : in STD_LOGIC_VECTOR(7 DOWNTO 0);
	  AddOut : out STD_LOGIC_VECTOR(7 DOWNTO 0));
END SomadorPC;

ARCHITECTURE behavior OF SomadorPC IS
BEGIN
	AddOut <= AddIn + AddInTwo;
END behavior;